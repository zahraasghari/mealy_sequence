library ieee ;
use ieee.std_logic_1164.all ;


entity mealy_sequence is

	port(
	
		clk : in std_logic ;
		input : in std_logic ;
		reset : in std_logic ;
		
		output : out std_logic 
	
	);

end mealy_sequence ;


architecture bhv of mealy_sequence is

	type state is (s0,s1,s2,s3,s4,s5) ;
	
	
	signal cs : state := s0 ;
	signal ns : state := s0 ;


begin

	process(clk ,reset )
	
	begin
	
		if reset = '1' then
		
			cs <= s0 ;
			
		elsif clk'event and clk = '1' then
		
			cs <= ns ;
			
		end if ;
	
	end process ;
	
	
	process(cs , input)
	
	begin
	
		case cs is
		
		when s0 =>
			
			if input = '1' then 
				ns <= s0;
				output <= '0' ;
			else 
				ns <= s1 ;
				output <= '0' ;
		
			end if ;
				
		when s1 =>
		
			if input = '1' then 
				ns <= s1 ;
				output <= '0' ;
			else 
				ns<= s2 ;
				output <= '0' ;
			end if ;
			
		when s2=>
			if input = '1' then 
				ns <= s3 ;
				output <= '0' ;
			else 
				ns <= s2 ;
				output <= '0' ;
			end if ;
       when s3 =>
			
			if input = '1' then 
				ns <= s4;
				output <= '0' ;
			else 
				ns <= s3 ;
				output <= '0' ;
		
			end if ;
				
		when s4 =>
		
			if input = '1' then 
				ns <= s4 ;
				output <= '0' ;
			else 
				ns <= s5 ;
				output <= '0' ;
			end if ;
			
		when s5=>
			if input = '1' then 
				ns <= s0 ;
				output <= '1' ;
			else 
				ns <= s2 ;
				output <= '0' ;
			end if ;
		end case ;
	
	end process ;






end bhv ;